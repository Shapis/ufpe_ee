LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE WORK.lcd_vhdl_package.ALL;
ENTITY lcd_logic IS
  PORT( 	clk      : IN  STD_LOGIC;  --clock principal			
			lcd_busy : IN  STD_LOGIC;  --feedback do controlador (1)ocupado/(0)disponível		
			--key		: IN 	STD_LOGIC_VECTOR(4 DOWNTO 1); --botões
			musica, autor : IN std_logic_vector (127 DOWNTO 0);
			lcd_e 	: OUT STD_LOGIC;  --retem os dados no controlador LCD
			lcd_bar	: OUT STD_LOGIC_VECTOR(9 DOWNTO 0)  --(9) rs (8) rw (7..0) dado char
		);
END lcd_logic;
ARCHITECTURE bhv OF lcd_logic IS
	--Registradores
	SIGNAL lcd_enable : STD_LOGIC;
	SIGNAL lcd_bus    : STD_LOGIC_VECTOR(9 DOWNTO 0);
	--Barramento de dados do display
	SIGNAL L1 : std_logic_vector (127 DOWNTO 0);
	SIGNAL L2 : std_logic_vector (127 DOWNTO 0);
BEGIN
	--atribuição contínua das saídas registradas
	lcd_e <= lcd_enable;
	lcd_bar <= lcd_bus; 
	
	--seleção do conteúdo através do key1
	L1 <= musica;
	L2 <= autor;

  --Sequenciamento do envio de cada caractere de L1 e L2
  PROCESS(clk)
    VARIABLE char  :  INTEGER RANGE 0 TO 34 := 0; --6 bits
  BEGIN
    IF rising_edge(clk) THEN
      IF (lcd_busy = '0' AND lcd_enable = '0') THEN
        lcd_enable <= '1'; --habilita o LCD
        IF (char < 34) THEN
          char := char + 1; --incrementa o estado
			ELSE char := 0; --reinicia o estado
        END IF;
        CASE char IS --verifica o estado atual
			 WHEN 0  => lcd_bus <= "00" & "10000000"; --inst. linha 1
          WHEN 1  => lcd_bus <= "10" & L1(127 DOWNTO 120); --prim. char da linha 1
          WHEN 2  => lcd_bus <= "10" & L1(119 DOWNTO 112);
          WHEN 3  => lcd_bus <= "10" & L1(111 DOWNTO 104);
          WHEN 4  => lcd_bus <= "10" & L1(103 DOWNTO 96);
          WHEN 5  => lcd_bus <= "10" & L1(95 DOWNTO 88);
          WHEN 6  => lcd_bus <= "10" & L1(87 DOWNTO 80);
          WHEN 7  => lcd_bus <= "10" & L1(79 DOWNTO 72);
          WHEN 8  => lcd_bus <= "10" & L1(71 DOWNTO 64);
          WHEN 9  => lcd_bus <= "10" & L1(63 DOWNTO 56);
			 WHEN 10 => lcd_bus <= "10" & L1(55 DOWNTO 48);
			 WHEN 11 => lcd_bus <= "10" & L1(47 DOWNTO 40);
			 WHEN 12 => lcd_bus <= "10" & L1(39 DOWNTO 32);
			 WHEN 13 => lcd_bus <= "10" & L1(31 DOWNTO 24);
			 WHEN 14 => lcd_bus <= "10" & L1(23 DOWNTO 16);
			 WHEN 15 => lcd_bus <= "10" & L1(15 DOWNTO 8);
			 WHEN 16 => lcd_bus <= "10" & L1(7 DOWNTO 0); --ult char da linha 1
			 WHEN 17 => lcd_bus <= "00" & "11000000"; --inst. linha 2
          WHEN 18 => lcd_bus <= "10" & L2(127 DOWNTO 120); --prim. char da linha 2
          WHEN 19 => lcd_bus <= "10" & L2(119 DOWNTO 112);
          WHEN 20 => lcd_bus <= "10" & L2(111 DOWNTO 104);
          WHEN 21 => lcd_bus <= "10" & L2(103 DOWNTO 96);
          WHEN 22 => lcd_bus <= "10" & L2(95 DOWNTO 88);
          WHEN 23 => lcd_bus <= "10" & L2(87 DOWNTO 80);
          WHEN 24 => lcd_bus <= "10" & L2(79 DOWNTO 72);
          WHEN 25 => lcd_bus <= "10" & L2(71 DOWNTO 64);
          WHEN 26 => lcd_bus <= "10" & L2(63 DOWNTO 56);
			 WHEN 27 => lcd_bus <= "10" & L2(55 DOWNTO 48);
			 WHEN 28 => lcd_bus <= "10" & L2(47 DOWNTO 40);
			 WHEN 29 => lcd_bus <= "10" & L2(39 DOWNTO 32);
			 WHEN 30 => lcd_bus <= "10" & L2(31 DOWNTO 24);
			 WHEN 31 => lcd_bus <= "10" & L2(23 DOWNTO 16);
			 WHEN 32 => lcd_bus <= "10" & L2(15 DOWNTO 8);
			 WHEN 33 => lcd_bus <= "10" & L2(7 DOWNTO 0);--ult. char da linha 2			 
          WHEN OTHERS => lcd_enable <= '0'; --desabilita o LCD
        END CASE;
      ELSE
        lcd_enable <= '0'; --desabilita o LCD
      END IF;
    END IF;
  END PROCESS;
END bhv;
